
// This module describes a adder,2 input adder (a + b)
// Make sure the widths are less than what is supported by the architecture
module ALU #(
                    parameter AWIDTH = 32,      // Width of adder's 1st input
                              BWIDTH = 32,      // Width of adder's 2nd input
                              PWIDTH = 32       // Output width
                   )
                   (
                    input [AWIDTH-1:0] a,  // adder input
                    input [BWIDTH-1:0] b,  // adder input
                    input sign,
                    input sub,
                    output [PWIDTH-1:0] p,  // Output
                    output overflow
                   );

  wire [PWIDTH-1:0] c;
  
  wire [BWIDTH-1:0] b_complement;

  assign b_complement = b ^ {32{sub}};

  assign p[ 0 ] = (a[ 0 ] & b[ 0 ] & sub) | (~a[ 0 ] & ~b[ 0 ] & sub) | (~a[ 0 ] & b[ 0 ] & ~sub) | (a[ 0 ] & ~b[ 0 ] & sub);
  assign c[ 0 ] = (a[ 0 ] & b[ 0 ]) | (~a[ 0 ] & b[ 0 ] & sub) | (a[ 0 ] & ~b[ 0 ] & sub);

  assign p[ 1 ] = (a[ 1 ] & b[ 1 ] & c[ 0 ]) | (~a[ 1 ] & ~b[ 1 ] & c[ 0 ]) | (~a[ 1 ] & b[ 1 ] & ~c[ 0 ]) | (a[ 1 ] & ~b[ 1 ] & ~c[ 0 ]);
  assign c[ 1 ] = (a[ 1 ] & b[ 1 ]) | (~a[ 1 ] & b[ 1 ] & c[ 0 ]) | (a[ 1 ] & ~b[ 1 ] & c[ 0 ]);

  assign p[ 2 ] = (a[ 2 ] & b[ 2 ] & c[ 1 ]) | (~a[ 2 ] & ~b[ 2 ] & c[ 1 ]) | (~a[ 2 ] & b[ 2 ] & ~c[ 1 ]) | (a[ 2 ] & ~b[ 2 ] & ~c[ 1 ]);
  assign c[ 2 ] = (a[ 2 ] & b[ 2 ]) | (~a[ 2 ] & b[ 2 ] & c[ 1 ]) | (a[ 2 ] & ~b[ 2 ] & c[ 1 ]);

  assign p[ 3 ] = (a[ 3 ] & b[ 3 ] & c[ 2 ]) | (~a[ 3 ] & ~b[ 3 ] & c[ 2 ]) | (~a[ 3 ] & b[ 3 ] & ~c[ 2 ]) | (a[ 3 ] & ~b[ 3 ] & ~c[ 2 ]);
  assign c[ 3 ] = (a[ 3 ] & b[ 3 ]) | (~a[ 3 ] & b[ 3 ] & c[ 2 ]) | (a[ 3 ] & ~b[ 3 ] & c[ 2 ]);

  assign p[ 4 ] = (a[ 4 ] & b[ 4 ] & c[ 3 ]) | (~a[ 4 ] & ~b[ 4 ] & c[ 3 ]) | (~a[ 4 ] & b[ 4 ] & ~c[ 3 ]) | (a[ 4 ] & ~b[ 4 ] & ~c[ 3 ]);
  assign c[ 4 ] = (a[ 4 ] & b[ 4 ]) | (~a[ 4 ] & b[ 4 ] & c[ 3 ]) | (a[ 4 ] & ~b[ 4 ] & c[ 3 ]);

  assign p[ 5 ] = (a[ 5 ] & b[ 5 ] & c[ 4 ]) | (~a[ 5 ] & ~b[ 5 ] & c[ 4 ]) | (~a[ 5 ] & b[ 5 ] & ~c[ 4 ]) | (a[ 5 ] & ~b[ 5 ] & ~c[ 4 ]);
  assign c[ 5 ] = (a[ 5 ] & b[ 5 ]) | (~a[ 5 ] & b[ 5 ] & c[ 4 ]) | (a[ 5 ] & ~b[ 5 ] & c[ 4 ]);

  assign p[ 6 ] = (a[ 6 ] & b[ 6 ] & c[ 5 ]) | (~a[ 6 ] & ~b[ 6 ] & c[ 5 ]) | (~a[ 6 ] & b[ 6 ] & ~c[ 5 ]) | (a[ 6 ] & ~b[ 6 ] & ~c[ 5 ]);
  assign c[ 6 ] = (a[ 6 ] & b[ 6 ]) | (~a[ 6 ] & b[ 6 ] & c[ 5 ]) | (a[ 6 ] & ~b[ 6 ] & c[ 5 ]);

  assign p[ 7 ] = (a[ 7 ] & b[ 7 ] & c[ 6 ]) | (~a[ 7 ] & ~b[ 7 ] & c[ 6 ]) | (~a[ 7 ] & b[ 7 ] & ~c[ 6 ]) | (a[ 7 ] & ~b[ 7 ] & ~c[ 6 ]);
  assign c[ 7 ] = (a[ 7 ] & b[ 7 ]) | (~a[ 7 ] & b[ 7 ] & c[ 6 ]) | (a[ 7 ] & ~b[ 7 ] & c[ 6 ]);

  assign p[ 8 ] = (a[ 8 ] & b[ 8 ] & c[ 7 ]) | (~a[ 8 ] & ~b[ 8 ] & c[ 7 ]) | (~a[ 8 ] & b[ 8 ] & ~c[ 7 ]) | (a[ 8 ] & ~b[ 8 ] & ~c[ 7 ]);
  assign c[ 8 ] = (a[ 8 ] & b[ 8 ]) | (~a[ 8 ] & b[ 8 ] & c[ 7 ]) | (a[ 8 ] & ~b[ 8 ] & c[ 7 ]);

  assign p[ 9 ] = (a[ 9 ] & b[ 9 ] & c[ 8 ]) | (~a[ 9 ] & ~b[ 9 ] & c[ 8 ]) | (~a[ 9 ] & b[ 9 ] & ~c[ 8 ]) | (a[ 9 ] & ~b[ 9 ] & ~c[ 8 ]);
  assign c[ 9 ] = (a[ 9 ] & b[ 9 ]) | (~a[ 9 ] & b[ 9 ] & c[ 8 ]) | (a[ 9 ] & ~b[ 9 ] & c[ 8 ]);

  assign p[ 10 ] = (a[ 10 ] & b[ 10 ] & c[ 9 ]) | (~a[ 10 ] & ~b[ 10 ] & c[ 9 ]) | (~a[ 10 ] & b[ 10 ] & ~c[ 9 ]) | (a[ 10 ] & ~b[ 10 ] & ~c[ 9 ]);
  assign c[ 10 ] = (a[ 10 ] & b[ 10 ]) | (~a[ 10 ] & b[ 10 ] & c[ 9 ]) | (a[ 10 ] & ~b[ 10 ] & c[ 9 ]);

  assign p[ 11 ] = (a[ 11 ] & b[ 11 ] & c[ 10 ]) | (~a[ 11 ] & ~b[ 11 ] & c[ 10 ]) | (~a[ 11 ] & b[ 11 ] & ~c[ 10 ]) | (a[ 11 ] & ~b[ 11 ] & ~c[ 10 ]);
  assign c[ 11 ] = (a[ 11 ] & b[ 11 ]) | (~a[ 11 ] & b[ 11 ] & c[ 10 ]) | (a[ 11 ] & ~b[ 11 ] & c[ 10 ]);

  assign p[ 12 ] = (a[ 12 ] & b[ 12 ] & c[ 11 ]) | (~a[ 12 ] & ~b[ 12 ] & c[ 11 ]) | (~a[ 12 ] & b[ 12 ] & ~c[ 11 ]) | (a[ 12 ] & ~b[ 12 ] & ~c[ 11 ]);
  assign c[ 12 ] = (a[ 12 ] & b[ 12 ]) | (~a[ 12 ] & b[ 12 ] & c[ 11 ]) | (a[ 12 ] & ~b[ 12 ] & c[ 11 ]);

  assign p[ 13 ] = (a[ 13 ] & b[ 13 ] & c[ 12 ]) | (~a[ 13 ] & ~b[ 13 ] & c[ 12 ]) | (~a[ 13 ] & b[ 13 ] & ~c[ 12 ]) | (a[ 13 ] & ~b[ 13 ] & ~c[ 12 ]);
  assign c[ 13 ] = (a[ 13 ] & b[ 13 ]) | (~a[ 13 ] & b[ 13 ] & c[ 12 ]) | (a[ 13 ] & ~b[ 13 ] & c[ 12 ]);

  assign p[ 14 ] = (a[ 14 ] & b[ 14 ] & c[ 13 ]) | (~a[ 14 ] & ~b[ 14 ] & c[ 13 ]) | (~a[ 14 ] & b[ 14 ] & ~c[ 13 ]) | (a[ 14 ] & ~b[ 14 ] & ~c[ 13 ]);
  assign c[ 14 ] = (a[ 14 ] & b[ 14 ]) | (~a[ 14 ] & b[ 14 ] & c[ 13 ]) | (a[ 14 ] & ~b[ 14 ] & c[ 13 ]);

  assign p[ 15 ] = (a[ 15 ] & b[ 15 ] & c[ 14 ]) | (~a[ 15 ] & ~b[ 15 ] & c[ 14 ]) | (~a[ 15 ] & b[ 15 ] & ~c[ 14 ]) | (a[ 15 ] & ~b[ 15 ] & ~c[ 14 ]);
  assign c[ 15 ] = (a[ 15 ] & b[ 15 ]) | (~a[ 15 ] & b[ 15 ] & c[ 14 ]) | (a[ 15 ] & ~b[ 15 ] & c[ 14 ]);

  assign p[ 16 ] = (a[ 16 ] & b[ 16 ] & c[ 15 ]) | (~a[ 16 ] & ~b[ 16 ] & c[ 15 ]) | (~a[ 16 ] & b[ 16 ] & ~c[ 15 ]) | (a[ 16 ] & ~b[ 16 ] & ~c[ 15 ]);
  assign c[ 16 ] = (a[ 16 ] & b[ 16 ]) | (~a[ 16 ] & b[ 16 ] & c[ 15 ]) | (a[ 16 ] & ~b[ 16 ] & c[ 15 ]);

  assign p[ 17 ] = (a[ 17 ] & b[ 17 ] & c[ 16 ]) | (~a[ 17 ] & ~b[ 17 ] & c[ 16 ]) | (~a[ 17 ] & b[ 17 ] & ~c[ 16 ]) | (a[ 17 ] & ~b[ 17 ] & ~c[ 16 ]);
  assign c[ 17 ] = (a[ 17 ] & b[ 17 ]) | (~a[ 17 ] & b[ 17 ] & c[ 16 ]) | (a[ 17 ] & ~b[ 17 ] & c[ 16 ]);

  assign p[ 18 ] = (a[ 18 ] & b[ 18 ] & c[ 17 ]) | (~a[ 18 ] & ~b[ 18 ] & c[ 17 ]) | (~a[ 18 ] & b[ 18 ] & ~c[ 17 ]) | (a[ 18 ] & ~b[ 18 ] & ~c[ 17 ]);
  assign c[ 18 ] = (a[ 18 ] & b[ 18 ]) | (~a[ 18 ] & b[ 18 ] & c[ 17 ]) | (a[ 18 ] & ~b[ 18 ] & c[ 17 ]);

  assign p[ 19 ] = (a[ 19 ] & b[ 19 ] & c[ 18 ]) | (~a[ 19 ] & ~b[ 19 ] & c[ 18 ]) | (~a[ 19 ] & b[ 19 ] & ~c[ 18 ]) | (a[ 19 ] & ~b[ 19 ] & ~c[ 18 ]);
  assign c[ 19 ] = (a[ 19 ] & b[ 19 ]) | (~a[ 19 ] & b[ 19 ] & c[ 18 ]) | (a[ 19 ] & ~b[ 19 ] & c[ 18 ]);

  assign p[ 20 ] = (a[ 20 ] & b[ 20 ] & c[ 19 ]) | (~a[ 20 ] & ~b[ 20 ] & c[ 19 ]) | (~a[ 20 ] & b[ 20 ] & ~c[ 19 ]) | (a[ 20 ] & ~b[ 20 ] & ~c[ 19 ]);
  assign c[ 20 ] = (a[ 20 ] & b[ 20 ]) | (~a[ 20 ] & b[ 20 ] & c[ 19 ]) | (a[ 20 ] & ~b[ 20 ] & c[ 19 ]);

  assign p[ 21 ] = (a[ 21 ] & b[ 21 ] & c[ 20 ]) | (~a[ 21 ] & ~b[ 21 ] & c[ 20 ]) | (~a[ 21 ] & b[ 21 ] & ~c[ 20 ]) | (a[ 21 ] & ~b[ 21 ] & ~c[ 20 ]);
  assign c[ 21 ] = (a[ 21 ] & b[ 21 ]) | (~a[ 21 ] & b[ 21 ] & c[ 20 ]) | (a[ 21 ] & ~b[ 21 ] & c[ 20 ]);

  assign p[ 22 ] = (a[ 22 ] & b[ 22 ] & c[ 21 ]) | (~a[ 22 ] & ~b[ 22 ] & c[ 21 ]) | (~a[ 22 ] & b[ 22 ] & ~c[ 21 ]) | (a[ 22 ] & ~b[ 22 ] & ~c[ 21 ]);
  assign c[ 22 ] = (a[ 22 ] & b[ 22 ]) | (~a[ 22 ] & b[ 22 ] & c[ 21 ]) | (a[ 22 ] & ~b[ 22 ] & c[ 21 ]);

  assign p[ 23 ] = (a[ 23 ] & b[ 23 ] & c[ 22 ]) | (~a[ 23 ] & ~b[ 23 ] & c[ 22 ]) | (~a[ 23 ] & b[ 23 ] & ~c[ 22 ]) | (a[ 23 ] & ~b[ 23 ] & ~c[ 22 ]);
  assign c[ 23 ] = (a[ 23 ] & b[ 23 ]) | (~a[ 23 ] & b[ 23 ] & c[ 22 ]) | (a[ 23 ] & ~b[ 23 ] & c[ 22 ]);

  assign p[ 24 ] = (a[ 24 ] & b[ 24 ] & c[ 23 ]) | (~a[ 24 ] & ~b[ 24 ] & c[ 23 ]) | (~a[ 24 ] & b[ 24 ] & ~c[ 23 ]) | (a[ 24 ] & ~b[ 24 ] & ~c[ 23 ]);
  assign c[ 24 ] = (a[ 24 ] & b[ 24 ]) | (~a[ 24 ] & b[ 24 ] & c[ 23 ]) | (a[ 24 ] & ~b[ 24 ] & c[ 23 ]);

  assign p[ 25 ] = (a[ 25 ] & b[ 25 ] & c[ 24 ]) | (~a[ 25 ] & ~b[ 25 ] & c[ 24 ]) | (~a[ 25 ] & b[ 25 ] & ~c[ 24 ]) | (a[ 25 ] & ~b[ 25 ] & ~c[ 24 ]);
  assign c[ 25 ] = (a[ 25 ] & b[ 25 ]) | (~a[ 25 ] & b[ 25 ] & c[ 24 ]) | (a[ 25 ] & ~b[ 25 ] & c[ 24 ]);

  assign p[ 26 ] = (a[ 26 ] & b[ 26 ] & c[ 25 ]) | (~a[ 26 ] & ~b[ 26 ] & c[ 25 ]) | (~a[ 26 ] & b[ 26 ] & ~c[ 25 ]) | (a[ 26 ] & ~b[ 26 ] & ~c[ 25 ]);
  assign c[ 26 ] = (a[ 26 ] & b[ 26 ]) | (~a[ 26 ] & b[ 26 ] & c[ 25 ]) | (a[ 26 ] & ~b[ 26 ] & c[ 25 ]);

  assign p[ 27 ] = (a[ 27 ] & b[ 27 ] & c[ 26 ]) | (~a[ 27 ] & ~b[ 27 ] & c[ 26 ]) | (~a[ 27 ] & b[ 27 ] & ~c[ 26 ]) | (a[ 27 ] & ~b[ 27 ] & ~c[ 26 ]);
  assign c[ 27 ] = (a[ 27 ] & b[ 27 ]) | (~a[ 27 ] & b[ 27 ] & c[ 26 ]) | (a[ 27 ] & ~b[ 27 ] & c[ 26 ]);

  assign p[ 28 ] = (a[ 28 ] & b[ 28 ] & c[ 27 ]) | (~a[ 28 ] & ~b[ 28 ] & c[ 27 ]) | (~a[ 28 ] & b[ 28 ] & ~c[ 27 ]) | (a[ 28 ] & ~b[ 28 ] & ~c[ 27 ]);
  assign c[ 28 ] = (a[ 28 ] & b[ 28 ]) | (~a[ 28 ] & b[ 28 ] & c[ 27 ]) | (a[ 28 ] & ~b[ 28 ] & c[ 27 ]);

  assign p[ 29 ] = (a[ 29 ] & b[ 29 ] & c[ 28 ]) | (~a[ 29 ] & ~b[ 29 ] & c[ 28 ]) | (~a[ 29 ] & b[ 29 ] & ~c[ 28 ]) | (a[ 29 ] & ~b[ 29 ] & ~c[ 28 ]);
  assign c[ 29 ] = (a[ 29 ] & b[ 29 ]) | (~a[ 29 ] & b[ 29 ] & c[ 28 ]) | (a[ 29 ] & ~b[ 29 ] & c[ 28 ]);

  assign p[ 30 ] = (a[ 30 ] & b[ 30 ] & c[ 29 ]) | (~a[ 30 ] & ~b[ 30 ] & c[ 29 ]) | (~a[ 30 ] & b[ 30 ] & ~c[ 29 ]) | (a[ 30 ] & ~b[ 30 ] & ~c[ 29 ]);
  assign c[ 30 ] = (a[ 30 ] & b[ 30 ]) | (~a[ 30 ] & b[ 30 ] & c[ 29 ]) | (a[ 30 ] & ~b[ 30 ] & c[ 29 ]);

  assign p[ 31 ] = (a[ 31 ] & b[ 31 ] & c[ 30 ]) | (~a[ 31 ] & ~b[ 31 ] & c[ 30 ]) | (~a[ 31 ] & b[ 31 ] & ~c[ 30 ]) | (a[ 31 ] & ~b[ 31 ] & ~c[ 30 ]);
  assign c[ 31 ] = (a[ 31 ] & b[ 31 ]) | (~a[ 31 ] & b[ 31 ] & c[ 30 ]) | (a[ 31 ] & ~b[ 31 ] & c[ 30 ]);

	assign overflow = sign ? (c[ 31 ] ^ c[ 30 ]) : (sub ^ c[ 31 ]); 		
  
endmodule